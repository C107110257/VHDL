-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"
-- CREATED		"Thu Nov 26 11:44:32 2020"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY sg IS 
	PORT
	(
		digit :  OUT  STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
END sg;

ARCHITECTURE bdf_type OF sg IS 

COMPONENT clk_src
	PORT(		 CLK : OUT STD_LOGIC;
		 RST : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT counter
	PORT(clk : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 digit : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;


BEGIN 



b2v_inst : clk_src
PORT MAP(		 CLK => SYNTHESIZED_WIRE_0,
		 RST => SYNTHESIZED_WIRE_1);


b2v_inst2 : counter
PORT MAP(clk => SYNTHESIZED_WIRE_0,
		 reset => SYNTHESIZED_WIRE_1,
		 digit => digit);


END bdf_type;