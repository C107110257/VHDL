LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
---------------------------------------
ENTITY ALU IS
	PORT( sel : IN STD_LOGIC_VECTOR(7 downto 0);
			square_output : OUT STD_LOGIC_VECTOR(7 downto 0);
			sawtooth_output : OUT STD_LOGIC_VECTOR(7 downto 0);
			triangle_output : OUT STD_LOGIC_VECTOR(7 downto 0);
			sine_output : OUT STD_LOGIC_VECTOR(7 downto 0));
END ALU;
---------------------------------------
ARCHITECTURE dataflow OF ALU IS
SIGNAL square, sawtooth, triangle, sine: STD_LOGIC_VECTOR(7 downto 0);
BEGIN
-----triangle unit:-----
	
	WITH sel(5 downto 0) SELECT
		triangle <= "00000001"  WHEN "000000",
						"00000010"  WHEN "000001",
						"00000011"  WHEN "000010",
						"00000100"  WHEN "000011",
						"00000101"  WHEN "000100",
						"00000110"  WHEN "000101",
						"00000111"  WHEN "000110",
						"00001000"  WHEN "000111",
						"00001001"  WHEN "001000",
						"00001010"  WHEN "001001",
						"00001011"  WHEN "001010",
						"00001100"  WHEN "001011",
						"00001101"  WHEN "001100",
						"00001110"  WHEN "001101",
						"00001111"  WHEN "001110",
						"00010000"  WHEN "001111",
						"00010001"  WHEN "010000",
						"00010010"  WHEN "010001",
						"00010011"  WHEN "010010",
						"00010100"  WHEN "010011",
						"00010101"  WHEN "010100",
						"00010110"  WHEN "010101",
						"00010111"  WHEN "010110",
						"00011000"  WHEN "010111",
						"00011001"  WHEN "011000",
						"00011010"  WHEN "011001",
						"00011011"  WHEN "011010",
						"00011100"  WHEN "011011",
						"00011101"  WHEN "011100",
						"00011110"  WHEN "011101",
						"00011111"  WHEN "011110",
						"00100000"  WHEN "011111",
						
						"00011111"  WHEN "100000",
						"00011110"  WHEN "100001",
						"00011101"  WHEN "100010",
						"00011100"  WHEN "100011",
						"00011011"  WHEN "100100",
						"00011010"  WHEN "100101",
						"00011001"  WHEN "100110",
						"00011000"  WHEN "100111",
						"00010111"  WHEN "101000",
						"00010110"  WHEN "101001",
						"00010101"  WHEN "101010",
						"00010100"  WHEN "101011",
						"00010011"  WHEN "101100",
						"00010010"  WHEN "101101",
						"00010001"  WHEN "101110",
						"00010000"  WHEN "101111",
						"00001111"  WHEN "110000",
						"00001110"  WHEN "110001",
						"00001101"  WHEN "110010",
						"00001100"  WHEN "110011",
						"00001011"  WHEN "110100",
						"00001010"  WHEN "110101",
						"00001001"  WHEN "110110",
						"00001000"  WHEN "110111",
						"00000111"  WHEN "111000",
						"00000110"  WHEN "111001",
						"00000101"  WHEN "111010",
						"00000100"  WHEN "111011",
						"00000011"  WHEN "111100",
						"00000010"  WHEN "111101",
						"00000001"  WHEN "111110",
						"00000000"  WHEN OTHERS;

-----sawtooth unit:-----
	WITH sel(5 downto 0) SELECT
		sawtooth <= "00000001"  WHEN "000000",
						"00000010"  WHEN "000001",
						"00000011"  WHEN "000010",
						"00000100"  WHEN "000011",
						"00000101"  WHEN "000100",
						"00000110"  WHEN "000101",
						"00000111"  WHEN "000110",
						"00001000"  WHEN "000111",
						"00001001"  WHEN "001000",
						"00001010"  WHEN "001001",
						"00001011"  WHEN "001010",
						"00001100"  WHEN "001011",
						"00001101"  WHEN "001100",
						"00001110"  WHEN "001101",
						"00001111"  WHEN "001110",
						"00010000"  WHEN "001111",
						"00010001"  WHEN "010000",
						"00010010"  WHEN "010001",
						"00010011"  WHEN "010010",
						"00010100"  WHEN "010011",
						"00010101"  WHEN "010100",
						"00010110"  WHEN "010101",
						"00010111"  WHEN "010110",
						"00011000"  WHEN "010111",
						"00011001"  WHEN "011000",
						"00011010"  WHEN "011001",
						"00011011"  WHEN "011010",
						"00011100"  WHEN "011011",
						"00011101"  WHEN "011100",
						"00011110"  WHEN "011101",
						"00011111"  WHEN "011110",
						"00100000"  WHEN "011111",
						
						"00100001"  WHEN "100000",
						"00100010"  WHEN "100001",
						"00100011"  WHEN "100010",
						"00100100"  WHEN "100011",
						"00100101"  WHEN "100100",
						"00100110"  WHEN "100101",
						"00100111"  WHEN "100110",
						"00101000"  WHEN "100111",
						"00101001"  WHEN "101000",
						"00101010"  WHEN "101001",
						"00101011"  WHEN "101010",
						"00101100"  WHEN "101011",
						"00101101"  WHEN "101100",
						"00101110"  WHEN "101101",
						"00101111"  WHEN "101110",
						"00110000"  WHEN "101111",
						"00110001"  WHEN "110000",
						"00110010"  WHEN "110001",
						"00110011"  WHEN "110010",
						"00110100"  WHEN "110011",
						"00110101"  WHEN "110100",
						"00110110"  WHEN "110101",
						"00110111"  WHEN "110110",
						"00111000"  WHEN "110111",
						"00111001"  WHEN "111000",
						"00111010"  WHEN "111001",
						"00111011"  WHEN "111010",
						"00111100"  WHEN "111011",
						"00111101"  WHEN "111100",
						"00111110"  WHEN "111101",
						"00111111"  WHEN "111110",
						"00000000"  WHEN OTHERS;
-----square unit:-----
	WITH sel(5 downto 0) SELECT
		square <= "00111111"  WHEN "000000",
						"00111111"  WHEN "000001",
						"00111111"  WHEN "000010",
						"00111111"  WHEN "000011",
						"00111111"  WHEN "000100",
						"00111111"  WHEN "000101",
						"00111111"  WHEN "000110",
						"00111111"  WHEN "000111",
						"00111111"  WHEN "001000",
						"00111111"  WHEN "001001",
						"00111111"  WHEN "001010",
						"00111111"  WHEN "001011",
						"00111111"  WHEN "001100",
						"00111111"  WHEN "001101",
						"00111111"  WHEN "001110",
						"00111111"  WHEN "001111",
						"00111111"  WHEN "010000",
						"00111111"  WHEN "010001",
						"00111111"  WHEN "010010",
						"00111111"  WHEN "010011",
						"00111111"  WHEN "010100",
						"00111111"  WHEN "010101",
						"00111111"  WHEN "010110",
						"00111111"  WHEN "010111",
						"00111111"  WHEN "011000",
						"00111111"  WHEN "011001",
						"00111111"  WHEN "011010",
						"00111111"  WHEN "011011",
						"00111111"  WHEN "011100",
						"00111111"  WHEN "011101",
						"00111111"  WHEN "011110",
						"00111111"  WHEN "011111",
						
						"00000000"  WHEN "100000",
						"00000000"  WHEN "100001",
						"00000000"  WHEN "100010",
						"00000000"  WHEN "100011",
						"00000000"  WHEN "100100",
						"00000000"  WHEN "100101",
						"00000000"  WHEN "100110",
						"00000000"  WHEN "100111",
						"00000000"  WHEN "101000",
						"00000000"  WHEN "101001",
						"00000000"  WHEN "101010",
						"00000000"  WHEN "101011",
						"00000000"  WHEN "101100",
						"00000000"  WHEN "101101",
						"00000000"  WHEN "101110",
						"00000000"  WHEN "101111",
						"00000000"  WHEN "110000",
						"00000000"  WHEN "110001",
						"00000000"  WHEN "110010",
						"00000000"  WHEN "110011",
						"00000000"  WHEN "110100",
						"00000000"  WHEN "110101",
						"00000000"  WHEN "110110",
						"00000000"  WHEN "110111",
						"00000000"  WHEN "111000",
						"00000000"  WHEN "111001",
						"00000000"  WHEN "111010",
						"00000000"  WHEN "111011",
						"00000000"  WHEN "111100",
						"00000000"  WHEN "111101",
						"00000000"  WHEN "111110",
						"00000000"  WHEN OTHERS;
-----sine unit:-----
	WITH sel(5 downto 0) SELECT
		sine <= 		"11111101"  WHEN "000000",
						"00000011"  WHEN "000001",
						"00000111"  WHEN "000010",
						"00001010"  WHEN "000011",
						"00001101"  WHEN "000100",
						"00010011"  WHEN "000101",
						"00011001"  WHEN "000110",
						"00011110"  WHEN "000111",
						"00100100"  WHEN "001000",
						"00101001"  WHEN "001001",
						"00101101"  WHEN "001010",
						"00110010"  WHEN "001011",
						"00110101"  WHEN "001100",
						"00111000"  WHEN "001101",
						"00111011"  WHEN "001110",
						"00111101"  WHEN "001111",
						"00111110"  WHEN "010000",
						"00111111"  WHEN "010001",
						"00111111"  WHEN "010010",
						"00111110"  WHEN "010011",
						"00111101"  WHEN "010100",
						"00111011"  WHEN "010101",
						"00111001"  WHEN "010110",
						"00110110"  WHEN "010111",
						"00110010"  WHEN "011000",
						"00101110"  WHEN "011001",
						"00101010"  WHEN "011010",
						"00100101"  WHEN "011011",
						"00100000"  WHEN "011100",
						"00011010"  WHEN "011101",
						"00010100"  WHEN "011110",
						"00001110"  WHEN "011111",
						
						"00000110"  WHEN "100000",
						"11111011"  WHEN "100001",
						"11110101"  WHEN "100010",
						"11101111"  WHEN "100011",
						"11101001"  WHEN "100100",
						"11100011"  WHEN "100101",
						"11011110"  WHEN "100110",
						"11011000"  WHEN "100111",
						"11010100"  WHEN "101000",
						"11001111"  WHEN "101001",
						"11001100"  WHEN "101010",
						"11001000"  WHEN "101011",
						"11000110"  WHEN "101100",
						"11000100"  WHEN "101101",
						"11000010"  WHEN "101110",
						"11000001"  WHEN "101111",
						"11000001"  WHEN "110000",
						"11000001"  WHEN "110001",
						"11000010"  WHEN "110010",
						"11000100"  WHEN "110011",
						"11000110"  WHEN "110100",
						"11001001"  WHEN "110101",
						"11001101"  WHEN "110110",
						"11010000"  WHEN "110111",
						"11010101"  WHEN "111000",
						"11011010"  WHEN "111001",
						"11011111"  WHEN "111010",
						"11100100"  WHEN "111011",
						"11101010"  WHEN "111100",
						"11110000"  WHEN "111101",
						"11110100"  WHEN "111110",
						"11111010"  WHEN OTHERS;

-----Mux:-----
	--WITH sel(7 downto 6) SELECT
		sawtooth_output <= sawtooth; --WHEN "00";
	--WITH sel(7 downto 6) SELECT
		triangle_output <= triangle; --WHEN "01";
	--WITH sel(7 downto 6) SELECT
		square_output <= square; --WHEN "10";
	--WITH sel(7 downto 6) SELECT
		sine_output <= sine; --WHEN "11";
END dataflow;

