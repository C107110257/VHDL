-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"
-- CREATED		"Thu Nov 26 11:50:04 2020"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY full_adder2 IS 
	PORT
	(
		cin :  IN  STD_LOGIC;
		a :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		b :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		s :  OUT  STD_LOGIC;
		cout :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END full_adder2;

ARCHITECTURE bdf_type OF full_adder2 IS 

COMPONENT full_adder
	PORT(a : IN STD_LOGIC;
		 b : IN STD_LOGIC;
		 cin : IN STD_LOGIC;
		 s : OUT STD_LOGIC;
		 cout : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;


BEGIN 



b2v_inst : full_adder
PORT MAP(a => a(0),
		 b => b(0),
		 cin => cin,
		 s => SYNTHESIZED_WIRE_0,
		 cout => cout(0));


b2v_inst1 : full_adder
PORT MAP(a => a(1),
		 b => b(1),
		 cin => SYNTHESIZED_WIRE_0,
		 s => s,
		 cout => cout(1));


END bdf_type;