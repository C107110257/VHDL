-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"
-- CREATED		"Thu Nov 05 11:33:42 2020"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY tb_top IS 
	PORT
	(
		y :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END tb_top;

ARCHITECTURE bdf_type OF tb_top IS 

COMPONENT counter
	PORT(CLK : IN STD_LOGIC;
		 RST : IN STD_LOGIC;
		 Y : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT clk_src
	PORT(		 CLK : OUT STD_LOGIC;
		 RST : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;


BEGIN 



b2v_inst : counter
PORT MAP(CLK => SYNTHESIZED_WIRE_0,
		 RST => SYNTHESIZED_WIRE_1,
		 Y => y);


b2v_inst2 : clk_src
PORT MAP(		 CLK => SYNTHESIZED_WIRE_0,
		 RST => SYNTHESIZED_WIRE_1);


END bdf_type;